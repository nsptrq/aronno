magic
tech sky130A
magscale 1 2
timestamp 1729321553
<< nwell >>
rect -290 -89 1394 977
<< nsubdiff >>
rect -254 907 -194 941
rect 1298 907 1358 941
rect -254 881 -220 907
rect -254 -19 -220 7
rect 1324 881 1358 907
rect 1324 -19 1358 7
rect -254 -53 -194 -19
rect 1298 -53 1358 -19
<< nsubdiffcont >>
rect -194 907 1298 941
rect -254 7 -220 881
rect 1324 7 1358 881
rect -194 -53 1298 -19
<< locali >>
rect -254 907 -194 941
rect 1298 907 1358 941
rect -254 881 -220 907
rect -254 -19 -220 7
rect 1324 881 1358 907
rect 1324 -19 1358 7
rect -254 -53 -194 -19
rect 1298 -53 1358 -19
<< viali >>
rect 1324 7 1358 66
<< metal1 >>
rect -163 973 -111 979
rect -111 924 575 970
rect -163 915 -111 921
rect -154 835 -32 869
rect -154 711 -120 835
rect -66 788 -32 835
rect 100 826 110 878
rect 178 826 188 878
rect 529 875 575 924
rect 370 829 734 875
rect 916 826 926 878
rect 994 826 1004 878
rect 1136 835 1258 869
rect 1136 788 1170 835
rect -72 776 88 788
rect -72 600 -18 776
rect 34 600 88 776
rect -72 588 88 600
rect 200 588 360 788
rect 472 776 632 788
rect 472 600 526 776
rect 578 600 632 776
rect 472 588 632 600
rect 744 588 904 788
rect 1016 776 1176 788
rect 1016 600 1070 776
rect 1122 600 1176 776
rect 1224 730 1258 835
rect 1016 588 1176 600
rect 261 463 299 588
rect 805 463 843 588
rect 261 425 843 463
rect 261 300 299 425
rect 805 300 843 425
rect -72 288 88 300
rect -154 53 -120 146
rect -72 112 -18 288
rect 34 112 88 288
rect -72 100 88 112
rect 200 100 360 300
rect 472 277 632 300
rect 472 112 526 277
rect 578 112 632 277
rect 472 100 632 112
rect 744 100 904 300
rect 1016 288 1176 300
rect 1016 112 1070 288
rect 1122 112 1176 288
rect 1016 100 1176 112
rect -66 53 -32 100
rect -154 19 -32 53
rect 100 10 110 62
rect 178 10 188 62
rect 370 13 734 59
rect 529 -36 575 13
rect 916 10 926 62
rect 994 10 1004 62
rect 1136 53 1170 100
rect 1224 53 1258 143
rect 1136 19 1258 53
rect 1318 66 1364 78
rect 1318 7 1324 66
rect 1358 7 1364 66
rect 1318 -5 1364 7
rect 1209 -36 1215 -33
rect 529 -82 1215 -36
rect 1209 -85 1215 -82
rect 1267 -85 1273 -33
<< via1 >>
rect -163 921 -111 973
rect 110 826 178 878
rect 926 826 994 878
rect -18 600 34 776
rect 526 600 578 776
rect 1070 600 1122 776
rect -18 112 34 288
rect 526 112 578 277
rect 1070 112 1122 288
rect 110 10 178 62
rect 926 10 994 62
rect 1215 -85 1267 -33
<< metal2 >>
rect -169 921 -163 973
rect -111 921 -105 973
rect 955 921 1264 923
rect -160 12 -114 921
rect 110 878 1264 921
rect 110 816 178 826
rect 994 877 1264 878
rect 926 816 994 826
rect -18 776 34 786
rect -18 470 34 600
rect 524 776 580 786
rect 524 590 580 600
rect 1070 776 1122 786
rect 1070 470 1122 600
rect -18 418 1122 470
rect -20 288 36 298
rect -20 102 36 112
rect 526 277 578 418
rect 526 102 578 112
rect 1068 288 1124 298
rect 1068 102 1124 112
rect 110 62 178 72
rect -160 10 110 12
rect 926 62 994 72
rect -160 -33 994 10
rect 1218 -27 1264 877
rect 1215 -33 1267 -27
rect -160 -34 178 -33
rect 1215 -91 1267 -85
<< via2 >>
rect 524 600 526 776
rect 526 600 578 776
rect 578 600 580 776
rect -20 112 -18 288
rect -18 112 34 288
rect 34 112 36 288
rect 1068 112 1070 288
rect 1070 112 1122 288
rect 1122 112 1124 288
<< metal3 >>
rect 514 776 590 781
rect 514 600 524 776
rect 580 600 590 776
rect 514 595 590 600
rect 522 474 582 595
rect -22 414 1126 474
rect -22 293 38 414
rect 1066 293 1126 414
rect -30 288 46 293
rect -30 112 -20 288
rect 36 112 46 288
rect -30 107 46 112
rect 1058 288 1134 293
rect 1058 112 1068 288
rect 1124 112 1134 288
rect 1058 107 1134 112
use sky130_fd_pr__pfet_01v8_BH5GQ5  sky130_fd_pr__pfet_01v8_BH5GQ5_0
timestamp 1729320448
transform 1 0 552 0 1 688
box -552 -200 552 200
use sky130_fd_pr__pfet_01v8_BH5GQ5  sky130_fd_pr__pfet_01v8_BH5GQ5_1
timestamp 1729320448
transform 1 0 552 0 1 200
box -552 -200 552 200
use sky130_fd_pr__pfet_01v8_LA8JHL  sky130_fd_pr__pfet_01v8_LA8JHL_0
timestamp 1729320448
transform 1 0 -93 0 1 164
box -109 -164 109 198
use sky130_fd_pr__pfet_01v8_LA8JHL  sky130_fd_pr__pfet_01v8_LA8JHL_1
timestamp 1729320448
transform 1 0 1197 0 1 164
box -109 -164 109 198
use sky130_fd_pr__pfet_01v8_MA8JHN  sky130_fd_pr__pfet_01v8_MA8JHN_0
timestamp 1729320448
transform 1 0 -93 0 1 724
box -109 -198 109 164
use sky130_fd_pr__pfet_01v8_MA8JHN  sky130_fd_pr__pfet_01v8_MA8JHN_1
timestamp 1729320448
transform 1 0 1197 0 1 724
box -109 -198 109 164
<< labels >>
flabel metal2 13 514 13 514 0 FreeSans 1600 0 0 0 VOUT
port 0 nsew
flabel viali 1345 33 1345 33 0 FreeSans 1600 0 0 0 VDD
port 1 nsew
flabel metal1 545 36 545 36 0 FreeSans 1600 0 0 0 VIP
port 2 nsew
flabel metal1 549 850 549 850 0 FreeSans 1600 0 0 0 VIN
port 3 nsew
flabel metal3 1098 358 1098 358 0 FreeSans 1600 0 0 0 D6
port 4 nsew
flabel metal1 279 341 279 341 0 FreeSans 1600 0 0 0 s67
port 5 nsew
<< end >>

magic
tech sky130A
magscale 1 2
timestamp 1729320448
<< nwell >>
rect -654 -973 654 973
<< pmos >>
rect -458 554 -358 754
rect -186 554 -86 754
rect 86 554 186 754
rect 358 554 458 754
rect -458 118 -358 318
rect -186 118 -86 318
rect 86 118 186 318
rect 358 118 458 318
rect -458 -318 -358 -118
rect -186 -318 -86 -118
rect 86 -318 186 -118
rect 358 -318 458 -118
rect -458 -754 -358 -554
rect -186 -754 -86 -554
rect 86 -754 186 -554
rect 358 -754 458 -554
<< pdiff >>
rect -516 742 -458 754
rect -516 566 -504 742
rect -470 566 -458 742
rect -516 554 -458 566
rect -358 742 -300 754
rect -358 566 -346 742
rect -312 566 -300 742
rect -358 554 -300 566
rect -244 742 -186 754
rect -244 566 -232 742
rect -198 566 -186 742
rect -244 554 -186 566
rect -86 742 -28 754
rect -86 566 -74 742
rect -40 566 -28 742
rect -86 554 -28 566
rect 28 742 86 754
rect 28 566 40 742
rect 74 566 86 742
rect 28 554 86 566
rect 186 742 244 754
rect 186 566 198 742
rect 232 566 244 742
rect 186 554 244 566
rect 300 742 358 754
rect 300 566 312 742
rect 346 566 358 742
rect 300 554 358 566
rect 458 742 516 754
rect 458 566 470 742
rect 504 566 516 742
rect 458 554 516 566
rect -516 306 -458 318
rect -516 130 -504 306
rect -470 130 -458 306
rect -516 118 -458 130
rect -358 306 -300 318
rect -358 130 -346 306
rect -312 130 -300 306
rect -358 118 -300 130
rect -244 306 -186 318
rect -244 130 -232 306
rect -198 130 -186 306
rect -244 118 -186 130
rect -86 306 -28 318
rect -86 130 -74 306
rect -40 130 -28 306
rect -86 118 -28 130
rect 28 306 86 318
rect 28 130 40 306
rect 74 130 86 306
rect 28 118 86 130
rect 186 306 244 318
rect 186 130 198 306
rect 232 130 244 306
rect 186 118 244 130
rect 300 306 358 318
rect 300 130 312 306
rect 346 130 358 306
rect 300 118 358 130
rect 458 306 516 318
rect 458 130 470 306
rect 504 130 516 306
rect 458 118 516 130
rect -516 -130 -458 -118
rect -516 -306 -504 -130
rect -470 -306 -458 -130
rect -516 -318 -458 -306
rect -358 -130 -300 -118
rect -358 -306 -346 -130
rect -312 -306 -300 -130
rect -358 -318 -300 -306
rect -244 -130 -186 -118
rect -244 -306 -232 -130
rect -198 -306 -186 -130
rect -244 -318 -186 -306
rect -86 -130 -28 -118
rect -86 -306 -74 -130
rect -40 -306 -28 -130
rect -86 -318 -28 -306
rect 28 -130 86 -118
rect 28 -306 40 -130
rect 74 -306 86 -130
rect 28 -318 86 -306
rect 186 -130 244 -118
rect 186 -306 198 -130
rect 232 -306 244 -130
rect 186 -318 244 -306
rect 300 -130 358 -118
rect 300 -306 312 -130
rect 346 -306 358 -130
rect 300 -318 358 -306
rect 458 -130 516 -118
rect 458 -306 470 -130
rect 504 -306 516 -130
rect 458 -318 516 -306
rect -516 -566 -458 -554
rect -516 -742 -504 -566
rect -470 -742 -458 -566
rect -516 -754 -458 -742
rect -358 -566 -300 -554
rect -358 -742 -346 -566
rect -312 -742 -300 -566
rect -358 -754 -300 -742
rect -244 -566 -186 -554
rect -244 -742 -232 -566
rect -198 -742 -186 -566
rect -244 -754 -186 -742
rect -86 -566 -28 -554
rect -86 -742 -74 -566
rect -40 -742 -28 -566
rect -86 -754 -28 -742
rect 28 -566 86 -554
rect 28 -742 40 -566
rect 74 -742 86 -566
rect 28 -754 86 -742
rect 186 -566 244 -554
rect 186 -742 198 -566
rect 232 -742 244 -566
rect 186 -754 244 -742
rect 300 -566 358 -554
rect 300 -742 312 -566
rect 346 -742 358 -566
rect 300 -754 358 -742
rect 458 -566 516 -554
rect 458 -742 470 -566
rect 504 -742 516 -566
rect 458 -754 516 -742
<< pdiffc >>
rect -504 566 -470 742
rect -346 566 -312 742
rect -232 566 -198 742
rect -74 566 -40 742
rect 40 566 74 742
rect 198 566 232 742
rect 312 566 346 742
rect 470 566 504 742
rect -504 130 -470 306
rect -346 130 -312 306
rect -232 130 -198 306
rect -74 130 -40 306
rect 40 130 74 306
rect 198 130 232 306
rect 312 130 346 306
rect 470 130 504 306
rect -504 -306 -470 -130
rect -346 -306 -312 -130
rect -232 -306 -198 -130
rect -74 -306 -40 -130
rect 40 -306 74 -130
rect 198 -306 232 -130
rect 312 -306 346 -130
rect 470 -306 504 -130
rect -504 -742 -470 -566
rect -346 -742 -312 -566
rect -232 -742 -198 -566
rect -74 -742 -40 -566
rect 40 -742 74 -566
rect 198 -742 232 -566
rect 312 -742 346 -566
rect 470 -742 504 -566
<< nsubdiff >>
rect -618 903 -522 937
rect 522 903 618 937
rect -618 841 -584 903
rect 584 841 618 903
rect -618 -903 -584 -841
rect 584 -903 618 -841
rect -618 -937 -522 -903
rect 522 -937 618 -903
<< nsubdiffcont >>
rect -522 903 522 937
rect -618 -841 -584 841
rect 584 -841 618 841
rect -522 -937 522 -903
<< poly >>
rect -458 835 -358 851
rect -458 801 -442 835
rect -374 801 -358 835
rect -458 754 -358 801
rect -186 835 -86 851
rect -186 801 -170 835
rect -102 801 -86 835
rect -186 754 -86 801
rect 86 835 186 851
rect 86 801 102 835
rect 170 801 186 835
rect 86 754 186 801
rect 358 835 458 851
rect 358 801 374 835
rect 442 801 458 835
rect 358 754 458 801
rect -458 507 -358 554
rect -458 473 -442 507
rect -374 473 -358 507
rect -458 457 -358 473
rect -186 507 -86 554
rect -186 473 -170 507
rect -102 473 -86 507
rect -186 457 -86 473
rect 86 507 186 554
rect 86 473 102 507
rect 170 473 186 507
rect 86 457 186 473
rect 358 507 458 554
rect 358 473 374 507
rect 442 473 458 507
rect 358 457 458 473
rect -458 399 -358 415
rect -458 365 -442 399
rect -374 365 -358 399
rect -458 318 -358 365
rect -186 399 -86 415
rect -186 365 -170 399
rect -102 365 -86 399
rect -186 318 -86 365
rect 86 399 186 415
rect 86 365 102 399
rect 170 365 186 399
rect 86 318 186 365
rect 358 399 458 415
rect 358 365 374 399
rect 442 365 458 399
rect 358 318 458 365
rect -458 71 -358 118
rect -458 37 -442 71
rect -374 37 -358 71
rect -458 21 -358 37
rect -186 71 -86 118
rect -186 37 -170 71
rect -102 37 -86 71
rect -186 21 -86 37
rect 86 71 186 118
rect 86 37 102 71
rect 170 37 186 71
rect 86 21 186 37
rect 358 71 458 118
rect 358 37 374 71
rect 442 37 458 71
rect 358 21 458 37
rect -458 -37 -358 -21
rect -458 -71 -442 -37
rect -374 -71 -358 -37
rect -458 -118 -358 -71
rect -186 -37 -86 -21
rect -186 -71 -170 -37
rect -102 -71 -86 -37
rect -186 -118 -86 -71
rect 86 -37 186 -21
rect 86 -71 102 -37
rect 170 -71 186 -37
rect 86 -118 186 -71
rect 358 -37 458 -21
rect 358 -71 374 -37
rect 442 -71 458 -37
rect 358 -118 458 -71
rect -458 -365 -358 -318
rect -458 -399 -442 -365
rect -374 -399 -358 -365
rect -458 -415 -358 -399
rect -186 -365 -86 -318
rect -186 -399 -170 -365
rect -102 -399 -86 -365
rect -186 -415 -86 -399
rect 86 -365 186 -318
rect 86 -399 102 -365
rect 170 -399 186 -365
rect 86 -415 186 -399
rect 358 -365 458 -318
rect 358 -399 374 -365
rect 442 -399 458 -365
rect 358 -415 458 -399
rect -458 -473 -358 -457
rect -458 -507 -442 -473
rect -374 -507 -358 -473
rect -458 -554 -358 -507
rect -186 -473 -86 -457
rect -186 -507 -170 -473
rect -102 -507 -86 -473
rect -186 -554 -86 -507
rect 86 -473 186 -457
rect 86 -507 102 -473
rect 170 -507 186 -473
rect 86 -554 186 -507
rect 358 -473 458 -457
rect 358 -507 374 -473
rect 442 -507 458 -473
rect 358 -554 458 -507
rect -458 -801 -358 -754
rect -458 -835 -442 -801
rect -374 -835 -358 -801
rect -458 -851 -358 -835
rect -186 -801 -86 -754
rect -186 -835 -170 -801
rect -102 -835 -86 -801
rect -186 -851 -86 -835
rect 86 -801 186 -754
rect 86 -835 102 -801
rect 170 -835 186 -801
rect 86 -851 186 -835
rect 358 -801 458 -754
rect 358 -835 374 -801
rect 442 -835 458 -801
rect 358 -851 458 -835
<< polycont >>
rect -442 801 -374 835
rect -170 801 -102 835
rect 102 801 170 835
rect 374 801 442 835
rect -442 473 -374 507
rect -170 473 -102 507
rect 102 473 170 507
rect 374 473 442 507
rect -442 365 -374 399
rect -170 365 -102 399
rect 102 365 170 399
rect 374 365 442 399
rect -442 37 -374 71
rect -170 37 -102 71
rect 102 37 170 71
rect 374 37 442 71
rect -442 -71 -374 -37
rect -170 -71 -102 -37
rect 102 -71 170 -37
rect 374 -71 442 -37
rect -442 -399 -374 -365
rect -170 -399 -102 -365
rect 102 -399 170 -365
rect 374 -399 442 -365
rect -442 -507 -374 -473
rect -170 -507 -102 -473
rect 102 -507 170 -473
rect 374 -507 442 -473
rect -442 -835 -374 -801
rect -170 -835 -102 -801
rect 102 -835 170 -801
rect 374 -835 442 -801
<< locali >>
rect -618 903 -522 937
rect 522 903 618 937
rect -618 841 -584 903
rect 584 841 618 903
rect -458 801 -442 835
rect -374 801 -358 835
rect -186 801 -170 835
rect -102 801 -86 835
rect 86 801 102 835
rect 170 801 186 835
rect 358 801 374 835
rect 442 801 458 835
rect -504 742 -470 758
rect -504 550 -470 566
rect -346 742 -312 758
rect -346 550 -312 566
rect -232 742 -198 758
rect -232 550 -198 566
rect -74 742 -40 758
rect -74 550 -40 566
rect 40 742 74 758
rect 40 550 74 566
rect 198 742 232 758
rect 198 550 232 566
rect 312 742 346 758
rect 312 550 346 566
rect 470 742 504 758
rect 470 550 504 566
rect -458 473 -442 507
rect -374 473 -358 507
rect -186 473 -170 507
rect -102 473 -86 507
rect 86 473 102 507
rect 170 473 186 507
rect 358 473 374 507
rect 442 473 458 507
rect -458 365 -442 399
rect -374 365 -358 399
rect -186 365 -170 399
rect -102 365 -86 399
rect 86 365 102 399
rect 170 365 186 399
rect 358 365 374 399
rect 442 365 458 399
rect -504 306 -470 322
rect -504 114 -470 130
rect -346 306 -312 322
rect -346 114 -312 130
rect -232 306 -198 322
rect -232 114 -198 130
rect -74 306 -40 322
rect -74 114 -40 130
rect 40 306 74 322
rect 40 114 74 130
rect 198 306 232 322
rect 198 114 232 130
rect 312 306 346 322
rect 312 114 346 130
rect 470 306 504 322
rect 470 114 504 130
rect -458 37 -442 71
rect -374 37 -358 71
rect -186 37 -170 71
rect -102 37 -86 71
rect 86 37 102 71
rect 170 37 186 71
rect 358 37 374 71
rect 442 37 458 71
rect -458 -71 -442 -37
rect -374 -71 -358 -37
rect -186 -71 -170 -37
rect -102 -71 -86 -37
rect 86 -71 102 -37
rect 170 -71 186 -37
rect 358 -71 374 -37
rect 442 -71 458 -37
rect -504 -130 -470 -114
rect -504 -322 -470 -306
rect -346 -130 -312 -114
rect -346 -322 -312 -306
rect -232 -130 -198 -114
rect -232 -322 -198 -306
rect -74 -130 -40 -114
rect -74 -322 -40 -306
rect 40 -130 74 -114
rect 40 -322 74 -306
rect 198 -130 232 -114
rect 198 -322 232 -306
rect 312 -130 346 -114
rect 312 -322 346 -306
rect 470 -130 504 -114
rect 470 -322 504 -306
rect -458 -399 -442 -365
rect -374 -399 -358 -365
rect -186 -399 -170 -365
rect -102 -399 -86 -365
rect 86 -399 102 -365
rect 170 -399 186 -365
rect 358 -399 374 -365
rect 442 -399 458 -365
rect -458 -507 -442 -473
rect -374 -507 -358 -473
rect -186 -507 -170 -473
rect -102 -507 -86 -473
rect 86 -507 102 -473
rect 170 -507 186 -473
rect 358 -507 374 -473
rect 442 -507 458 -473
rect -504 -566 -470 -550
rect -504 -758 -470 -742
rect -346 -566 -312 -550
rect -346 -758 -312 -742
rect -232 -566 -198 -550
rect -232 -758 -198 -742
rect -74 -566 -40 -550
rect -74 -758 -40 -742
rect 40 -566 74 -550
rect 40 -758 74 -742
rect 198 -566 232 -550
rect 198 -758 232 -742
rect 312 -566 346 -550
rect 312 -758 346 -742
rect 470 -566 504 -550
rect 470 -758 504 -742
rect -458 -835 -442 -801
rect -374 -835 -358 -801
rect -186 -835 -170 -801
rect -102 -835 -86 -801
rect 86 -835 102 -801
rect 170 -835 186 -801
rect 358 -835 374 -801
rect 442 -835 458 -801
rect -618 -903 -584 -841
rect 584 -903 618 -841
rect -618 -937 -522 -903
rect 522 -937 618 -903
<< viali >>
rect -442 801 -374 835
rect -170 801 -102 835
rect 102 801 170 835
rect 374 801 442 835
rect -504 566 -470 742
rect -346 566 -312 742
rect -232 566 -198 742
rect -74 566 -40 742
rect 40 566 74 742
rect 198 566 232 742
rect 312 566 346 742
rect 470 566 504 742
rect -442 473 -374 507
rect -170 473 -102 507
rect 102 473 170 507
rect 374 473 442 507
rect -442 365 -374 399
rect -170 365 -102 399
rect 102 365 170 399
rect 374 365 442 399
rect -504 130 -470 306
rect -346 130 -312 306
rect -232 130 -198 306
rect -74 130 -40 306
rect 40 130 74 306
rect 198 130 232 306
rect 312 130 346 306
rect 470 130 504 306
rect -442 37 -374 71
rect -170 37 -102 71
rect 102 37 170 71
rect 374 37 442 71
rect -442 -71 -374 -37
rect -170 -71 -102 -37
rect 102 -71 170 -37
rect 374 -71 442 -37
rect -504 -306 -470 -130
rect -346 -306 -312 -130
rect -232 -306 -198 -130
rect -74 -306 -40 -130
rect 40 -306 74 -130
rect 198 -306 232 -130
rect 312 -306 346 -130
rect 470 -306 504 -130
rect -442 -399 -374 -365
rect -170 -399 -102 -365
rect 102 -399 170 -365
rect 374 -399 442 -365
rect -442 -507 -374 -473
rect -170 -507 -102 -473
rect 102 -507 170 -473
rect 374 -507 442 -473
rect -504 -742 -470 -566
rect -346 -742 -312 -566
rect -232 -742 -198 -566
rect -74 -742 -40 -566
rect 40 -742 74 -566
rect 198 -742 232 -566
rect 312 -742 346 -566
rect 470 -742 504 -566
rect -442 -835 -374 -801
rect -170 -835 -102 -801
rect 102 -835 170 -801
rect 374 -835 442 -801
<< metal1 >>
rect -454 835 -362 841
rect -454 801 -442 835
rect -374 801 -362 835
rect -454 795 -362 801
rect -182 835 -90 841
rect -182 801 -170 835
rect -102 801 -90 835
rect -182 795 -90 801
rect 90 835 182 841
rect 90 801 102 835
rect 170 801 182 835
rect 90 795 182 801
rect 362 835 454 841
rect 362 801 374 835
rect 442 801 454 835
rect 362 795 454 801
rect -510 742 -464 754
rect -510 566 -504 742
rect -470 566 -464 742
rect -510 554 -464 566
rect -352 742 -306 754
rect -352 566 -346 742
rect -312 566 -306 742
rect -352 554 -306 566
rect -238 742 -192 754
rect -238 566 -232 742
rect -198 566 -192 742
rect -238 554 -192 566
rect -80 742 -34 754
rect -80 566 -74 742
rect -40 566 -34 742
rect -80 554 -34 566
rect 34 742 80 754
rect 34 566 40 742
rect 74 566 80 742
rect 34 554 80 566
rect 192 742 238 754
rect 192 566 198 742
rect 232 566 238 742
rect 192 554 238 566
rect 306 742 352 754
rect 306 566 312 742
rect 346 566 352 742
rect 306 554 352 566
rect 464 742 510 754
rect 464 566 470 742
rect 504 566 510 742
rect 464 554 510 566
rect -454 507 -362 513
rect -454 473 -442 507
rect -374 473 -362 507
rect -454 467 -362 473
rect -182 507 -90 513
rect -182 473 -170 507
rect -102 473 -90 507
rect -182 467 -90 473
rect 90 507 182 513
rect 90 473 102 507
rect 170 473 182 507
rect 90 467 182 473
rect 362 507 454 513
rect 362 473 374 507
rect 442 473 454 507
rect 362 467 454 473
rect -454 399 -362 405
rect -454 365 -442 399
rect -374 365 -362 399
rect -454 359 -362 365
rect -182 399 -90 405
rect -182 365 -170 399
rect -102 365 -90 399
rect -182 359 -90 365
rect 90 399 182 405
rect 90 365 102 399
rect 170 365 182 399
rect 90 359 182 365
rect 362 399 454 405
rect 362 365 374 399
rect 442 365 454 399
rect 362 359 454 365
rect -510 306 -464 318
rect -510 130 -504 306
rect -470 130 -464 306
rect -510 118 -464 130
rect -352 306 -306 318
rect -352 130 -346 306
rect -312 130 -306 306
rect -352 118 -306 130
rect -238 306 -192 318
rect -238 130 -232 306
rect -198 130 -192 306
rect -238 118 -192 130
rect -80 306 -34 318
rect -80 130 -74 306
rect -40 130 -34 306
rect -80 118 -34 130
rect 34 306 80 318
rect 34 130 40 306
rect 74 130 80 306
rect 34 118 80 130
rect 192 306 238 318
rect 192 130 198 306
rect 232 130 238 306
rect 192 118 238 130
rect 306 306 352 318
rect 306 130 312 306
rect 346 130 352 306
rect 306 118 352 130
rect 464 306 510 318
rect 464 130 470 306
rect 504 130 510 306
rect 464 118 510 130
rect -454 71 -362 77
rect -454 37 -442 71
rect -374 37 -362 71
rect -454 31 -362 37
rect -182 71 -90 77
rect -182 37 -170 71
rect -102 37 -90 71
rect -182 31 -90 37
rect 90 71 182 77
rect 90 37 102 71
rect 170 37 182 71
rect 90 31 182 37
rect 362 71 454 77
rect 362 37 374 71
rect 442 37 454 71
rect 362 31 454 37
rect -454 -37 -362 -31
rect -454 -71 -442 -37
rect -374 -71 -362 -37
rect -454 -77 -362 -71
rect -182 -37 -90 -31
rect -182 -71 -170 -37
rect -102 -71 -90 -37
rect -182 -77 -90 -71
rect 90 -37 182 -31
rect 90 -71 102 -37
rect 170 -71 182 -37
rect 90 -77 182 -71
rect 362 -37 454 -31
rect 362 -71 374 -37
rect 442 -71 454 -37
rect 362 -77 454 -71
rect -510 -130 -464 -118
rect -510 -306 -504 -130
rect -470 -306 -464 -130
rect -510 -318 -464 -306
rect -352 -130 -306 -118
rect -352 -306 -346 -130
rect -312 -306 -306 -130
rect -352 -318 -306 -306
rect -238 -130 -192 -118
rect -238 -306 -232 -130
rect -198 -306 -192 -130
rect -238 -318 -192 -306
rect -80 -130 -34 -118
rect -80 -306 -74 -130
rect -40 -306 -34 -130
rect -80 -318 -34 -306
rect 34 -130 80 -118
rect 34 -306 40 -130
rect 74 -306 80 -130
rect 34 -318 80 -306
rect 192 -130 238 -118
rect 192 -306 198 -130
rect 232 -306 238 -130
rect 192 -318 238 -306
rect 306 -130 352 -118
rect 306 -306 312 -130
rect 346 -306 352 -130
rect 306 -318 352 -306
rect 464 -130 510 -118
rect 464 -306 470 -130
rect 504 -306 510 -130
rect 464 -318 510 -306
rect -454 -365 -362 -359
rect -454 -399 -442 -365
rect -374 -399 -362 -365
rect -454 -405 -362 -399
rect -182 -365 -90 -359
rect -182 -399 -170 -365
rect -102 -399 -90 -365
rect -182 -405 -90 -399
rect 90 -365 182 -359
rect 90 -399 102 -365
rect 170 -399 182 -365
rect 90 -405 182 -399
rect 362 -365 454 -359
rect 362 -399 374 -365
rect 442 -399 454 -365
rect 362 -405 454 -399
rect -454 -473 -362 -467
rect -454 -507 -442 -473
rect -374 -507 -362 -473
rect -454 -513 -362 -507
rect -182 -473 -90 -467
rect -182 -507 -170 -473
rect -102 -507 -90 -473
rect -182 -513 -90 -507
rect 90 -473 182 -467
rect 90 -507 102 -473
rect 170 -507 182 -473
rect 90 -513 182 -507
rect 362 -473 454 -467
rect 362 -507 374 -473
rect 442 -507 454 -473
rect 362 -513 454 -507
rect -510 -566 -464 -554
rect -510 -742 -504 -566
rect -470 -742 -464 -566
rect -510 -754 -464 -742
rect -352 -566 -306 -554
rect -352 -742 -346 -566
rect -312 -742 -306 -566
rect -352 -754 -306 -742
rect -238 -566 -192 -554
rect -238 -742 -232 -566
rect -198 -742 -192 -566
rect -238 -754 -192 -742
rect -80 -566 -34 -554
rect -80 -742 -74 -566
rect -40 -742 -34 -566
rect -80 -754 -34 -742
rect 34 -566 80 -554
rect 34 -742 40 -566
rect 74 -742 80 -566
rect 34 -754 80 -742
rect 192 -566 238 -554
rect 192 -742 198 -566
rect 232 -742 238 -566
rect 192 -754 238 -742
rect 306 -566 352 -554
rect 306 -742 312 -566
rect 346 -742 352 -566
rect 306 -754 352 -742
rect 464 -566 510 -554
rect 464 -742 470 -566
rect 504 -742 510 -566
rect 464 -754 510 -742
rect -454 -801 -362 -795
rect -454 -835 -442 -801
rect -374 -835 -362 -801
rect -454 -841 -362 -835
rect -182 -801 -90 -795
rect -182 -835 -170 -801
rect -102 -835 -90 -801
rect -182 -841 -90 -835
rect 90 -801 182 -795
rect 90 -835 102 -801
rect 170 -835 182 -801
rect 90 -841 182 -835
rect 362 -801 454 -795
rect 362 -835 374 -801
rect 442 -835 454 -801
rect 362 -841 454 -835
<< properties >>
string FIXED_BBOX -601 -920 601 920
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 1 l 0.5 m 4 nf 4 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 0 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>

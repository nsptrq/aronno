magic
tech sky130A
magscale 1 2
timestamp 1729243325
<< pwell >>
rect -353 -785 1023 644
<< psubdiff >>
rect -290 577 -230 611
rect 918 577 978 611
rect -290 551 -256 577
rect 944 551 978 577
rect -290 -731 -256 -705
rect 944 -731 978 -705
rect -290 -765 -230 -731
rect 918 -765 978 -731
<< psubdiffcont >>
rect -230 577 918 611
rect -290 -705 -256 551
rect 944 -705 978 551
rect -230 -765 918 -731
<< poly >>
rect 58 -129 630 -20
<< locali >>
rect -290 577 -230 611
rect 918 577 978 611
rect -290 551 -256 577
rect 944 551 978 577
rect -102 458 -68 530
rect 756 458 790 530
rect 756 -684 790 -552
rect -290 -731 -256 -705
rect 944 -731 978 -705
rect -290 -765 -230 -731
rect 918 -765 978 -731
<< viali >>
rect 270 577 304 611
<< metal1 >>
rect 258 611 316 617
rect 258 577 270 611
rect 304 577 316 611
rect 258 571 316 577
rect -108 458 -62 530
rect -196 58 -62 458
rect 270 446 304 571
rect 750 458 796 530
rect 6 58 52 98
rect 251 70 261 446
rect 313 70 323 446
rect 365 70 375 446
rect 427 70 437 446
rect -108 26 52 58
rect 636 58 682 87
rect 750 58 884 458
rect -108 12 108 26
rect 6 -20 108 12
rect 636 12 796 58
rect 636 -54 682 12
rect 6 -100 682 -54
rect 6 -166 52 -100
rect -108 -212 52 -166
rect 595 -167 682 -134
rect 595 -180 796 -167
rect -196 -612 -62 -212
rect 6 -214 52 -212
rect 636 -212 796 -180
rect 636 -213 884 -212
rect 251 -600 261 -224
rect 313 -600 323 -224
rect 365 -600 375 -224
rect 427 -600 437 -224
rect 750 -612 884 -213
rect -108 -684 -62 -612
rect 756 -684 790 -612
<< via1 >>
rect 261 70 313 446
rect 375 70 427 446
rect 261 -600 313 -224
rect 375 -600 427 -224
<< metal2 >>
rect 261 446 313 456
rect 261 -50 313 70
rect 373 446 429 456
rect 373 60 429 70
rect 261 -102 427 -50
rect 259 -224 315 -214
rect 259 -610 315 -600
rect 375 -224 427 -102
rect 375 -610 427 -600
<< via2 >>
rect 373 70 375 446
rect 375 70 427 446
rect 427 70 429 446
rect 259 -600 261 -224
rect 261 -600 313 -224
rect 313 -600 315 -224
<< metal3 >>
rect 363 446 439 451
rect 363 70 373 446
rect 429 70 439 446
rect 363 65 439 70
rect 371 -46 431 65
rect 257 -106 431 -46
rect 257 -219 317 -106
rect 249 -224 325 -219
rect 249 -600 259 -224
rect 315 -600 325 -224
rect 249 -605 325 -600
use sky130_fd_pr__nfet_01v8_7CP4KT  sky130_fd_pr__nfet_01v8_7CP4KT_0
timestamp 1729238886
transform 1 0 -129 0 1 289
box -73 -257 73 257
use sky130_fd_pr__nfet_01v8_7CP4KT  sky130_fd_pr__nfet_01v8_7CP4KT_1
timestamp 1729238886
transform 1 0 817 0 1 289
box -73 -257 73 257
use sky130_fd_pr__nfet_01v8_7CYQ2Z  sky130_fd_pr__nfet_01v8_7CYQ2Z_0
timestamp 1729238886
transform 1 0 -129 0 1 -443
box -73 -257 73 257
use sky130_fd_pr__nfet_01v8_7CYQ2Z  sky130_fd_pr__nfet_01v8_7CYQ2Z_1
timestamp 1729238886
transform 1 0 817 0 1 -443
box -73 -257 73 257
use sky130_fd_pr__nfet_01v8_8UMB6F  sky130_fd_pr__nfet_01v8_8UMB6F_0
timestamp 1729238886
transform 1 0 344 0 1 -412
box -344 -288 344 288
use sky130_fd_pr__nfet_01v8_8UMB6F  sky130_fd_pr__nfet_01v8_8UMB6F_1
timestamp 1729238886
transform 1 0 344 0 1 258
box -344 -288 344 288
<< labels >>
flabel metal1 290 566 290 566 0 FreeSans 1600 0 0 0 GND
port 0 nsew
flabel metal1 -110 124 -110 124 0 FreeSans 1600 0 0 0 D3
port 1 nsew
flabel metal1 -106 -340 -106 -340 0 FreeSans 1600 0 0 0 D4
port 2 nsew
flabel metal3 276 -210 276 -210 0 FreeSans 1600 0 0 0 RS
port 3 nsew
<< end >>

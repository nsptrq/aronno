** sch_path: /home/nsptrq/newproject/ringosci/ringosci.sch
**.subckt ringosci vdd out gnd
*.iopin out
*.iopin vdd
*.iopin gnd
x1 vdd out net1 gnd inverter
x2 vdd net1 net2 gnd inverter
x3 vdd net2 out gnd inverter
**.ends

* expanding   symbol:  /home/nsptrq/newproject/inverter/inverter.sym # of pins=4
** sym_path: /home/nsptrq/newproject/inverter/inverter.sym
** sch_path: /home/nsptrq/newproject/inverter/inverter.sch
.subckt inverter vdd in out gnd
*.ipin vdd
*.ipin in
*.ipin gnd
*.opin out
XM1 out in gnd gnd sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM2 out in vdd vdd sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
.ends

.end

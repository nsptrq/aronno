magic
tech sky130A
magscale 1 2
timestamp 1729416081
<< nwell >>
rect -725 3938 255 4202
rect 1048 4076 1057 4087
rect 1042 3238 1062 3284
rect -725 842 273 1095
<< viali >>
rect 203 3296 237 3355
rect 291 3296 325 3355
rect 1027 2205 1061 2239
<< metal1 >>
rect 1048 4076 1057 4087
rect 1609 3722 1615 3774
rect 1667 3722 1964 3774
rect 2016 3722 2026 3774
rect 197 3355 243 3367
rect 285 3355 331 3367
rect 197 3296 203 3355
rect 237 3296 291 3355
rect 325 3296 331 3355
rect 197 3284 243 3296
rect 285 3284 331 3296
rect 808 3167 842 3388
rect 1042 3238 1062 3284
rect 1859 3232 1917 3281
rect 385 3133 842 3167
rect -4 2684 6 3060
rect 58 2684 68 3060
rect 385 2594 419 3133
rect 596 2731 656 2737
rect 656 2684 848 2718
rect 596 2665 656 2671
rect 370 2542 376 2594
rect 428 2542 434 2594
rect 4 2420 10 2472
rect 62 2469 68 2472
rect 62 2423 446 2469
rect 62 2420 68 2423
rect 400 1686 446 2423
rect 1027 2245 1061 2327
rect 1015 2239 1073 2245
rect 1015 2205 1027 2239
rect 1061 2205 1073 2239
rect 1015 2199 1073 2205
rect 400 1640 862 1686
rect 806 1475 871 1481
rect 806 1404 871 1410
<< via1 >>
rect 1615 3722 1667 3774
rect 1964 3722 2016 3774
rect 6 2684 58 3060
rect 596 2671 656 2731
rect 376 2542 428 2594
rect 10 2420 62 2472
rect 806 1410 871 1475
<< metal2 >>
rect 1615 3774 1667 3780
rect 1615 3716 1667 3722
rect 1962 3776 2018 3786
rect 1962 3710 2018 3720
rect 4 3060 60 3070
rect 525 2731 581 2738
rect 4 2674 60 2684
rect 523 2729 596 2731
rect 523 2673 525 2729
rect 581 2673 596 2729
rect 523 2671 596 2673
rect 656 2671 662 2731
rect 1948 2715 1957 2718
rect 525 2664 581 2671
rect 1674 2656 1957 2715
rect 1948 2652 1957 2656
rect 2023 2652 2032 2718
rect 376 2594 428 2600
rect 103 2551 376 2585
rect 376 2536 428 2542
rect 10 2472 62 2478
rect 10 2414 62 2420
rect 300 1475 356 1479
rect 296 1470 806 1475
rect 296 1414 300 1470
rect 356 1414 806 1470
rect 296 1410 806 1414
rect 871 1410 877 1475
rect 300 1405 356 1410
<< via2 >>
rect 1962 3774 2018 3776
rect 1962 3722 1964 3774
rect 1964 3722 2016 3774
rect 2016 3722 2018 3774
rect 1962 3720 2018 3722
rect 4 2684 6 3060
rect 6 2684 58 3060
rect 58 2684 60 3060
rect 525 2673 581 2729
rect 1957 2652 2023 2718
rect 300 1414 356 1470
<< metal3 >>
rect 1952 3776 2028 3781
rect 1952 3720 1962 3776
rect 2018 3720 2028 3776
rect -6 3060 70 3065
rect -6 2684 4 3060
rect 60 2750 70 3060
rect 60 2685 360 2750
rect 523 2734 583 3387
rect 60 2684 70 2685
rect -6 2679 70 2684
rect 295 1475 360 2685
rect 520 2729 586 2734
rect 520 2673 525 2729
rect 581 2673 586 2729
rect 520 2668 586 2673
rect 1952 2718 2028 3720
rect 1952 2652 1957 2718
rect 2023 2652 2028 2718
rect 1952 2647 2028 2652
rect 1302 1628 1338 1668
rect 295 1470 361 1475
rect 295 1414 300 1470
rect 356 1414 361 1470
rect 295 1409 361 1414
use nmoscs  nmoscs_0
timestamp 1729243325
transform 1 0 924 0 1 1628
box -353 -785 1023 644
use nmosout  nmosout_0
timestamp 1729332766
transform 1 0 797 0 1 2358
box -176 -77 1106 757
use pmoscs  pmoscs_0
timestamp 1729225119
transform 1 0 -559 0 1 1202
box -166 -107 832 2753
use pmosout  pmosout_0
timestamp 1729321553
transform 1 0 545 0 1 3225
box -290 -91 1394 979
<< labels >>
flabel metal3 1320 1648 1320 1648 0 FreeSans 1600 0 0 0 rs
port 0 nsew
flabel metal1 1043 2258 1043 2258 0 FreeSans 1600 0 0 0 gnd
port 1 nsew
flabel metal3 1980 2909 1980 2909 0 FreeSans 1600 0 0 0 vout
port 2 nsew
flabel metal1 1914 3241 1914 3241 0 FreeSans 1600 0 0 0 vdd
port 3 nsew
flabel metal1 1055 3262 1055 3262 0 FreeSans 1600 0 0 0 vip
port 4 nsew
flabel metal1 1053 4082 1053 4082 0 FreeSans 1600 0 0 0 vin
port 5 nsew
<< end >>

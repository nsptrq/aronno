magic
tech sky130A
magscale 1 2
timestamp 1729423519
use sky130_fd_pr__nfet_01v8_M9466H  sky130_fd_pr__nfet_01v8_M9466H_0
timestamp 1729423519
transform 1 0 835 0 1 357
box -296 -410 296 410
use sky130_fd_pr__pfet_01v8_LXK9WL  sky130_fd_pr__pfet_01v8_LXK9WL_0
timestamp 1729423519
transform 1 0 243 0 1 366
box -296 -419 296 419
<< end >>

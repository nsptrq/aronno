magic
tech sky130A
magscale 1 2
timestamp 1729225119
<< nwell >>
rect -166 -107 832 2753
<< nsubdiff >>
rect -130 2683 -70 2717
rect 736 2683 796 2717
rect -130 2657 -96 2683
rect 762 2657 796 2683
rect -130 -37 -96 -11
rect 762 -37 796 -11
rect -130 -71 -70 -37
rect 736 -71 796 -37
<< nsubdiffcont >>
rect -70 2683 736 2717
rect -130 -11 -96 2657
rect 762 -11 796 2657
rect -70 -71 736 -37
<< poly >>
rect -46 2645 46 2661
rect -46 2611 -30 2645
rect 4 2611 46 2645
rect -46 2595 46 2611
rect 16 2564 46 2595
rect 620 2645 712 2661
rect 620 2611 662 2645
rect 696 2611 712 2645
rect 620 2595 712 2611
rect 620 2588 650 2595
rect -46 1951 46 1967
rect 104 1965 304 2069
rect -46 1917 -30 1951
rect 4 1917 46 1951
rect -46 1901 46 1917
rect 16 1870 46 1901
rect 620 1951 712 1967
rect 620 1917 662 1951
rect 696 1917 712 1951
rect 620 1901 712 1917
rect 620 1870 650 1901
rect 104 1270 562 1379
rect 16 745 46 776
rect -46 729 46 745
rect -46 695 -30 729
rect 4 695 46 729
rect -46 679 46 695
rect 620 745 650 776
rect 620 729 712 745
rect 620 695 662 729
rect 696 695 712 729
rect 362 574 562 684
rect 620 679 712 695
rect 16 51 46 82
rect -46 35 46 51
rect -46 1 -30 35
rect 4 1 46 35
rect -46 -15 46 1
rect 620 51 650 82
rect 620 35 712 51
rect 620 1 662 35
rect 696 1 712 35
rect 620 -15 712 1
<< polycont >>
rect -30 2611 4 2645
rect 662 2611 696 2645
rect -30 1917 4 1951
rect 662 1917 696 1951
rect -30 695 4 729
rect 662 695 696 729
rect -30 1 4 35
rect 662 1 696 35
<< locali >>
rect -130 2683 -70 2717
rect 736 2683 796 2717
rect -130 2657 -96 2683
rect 762 2657 796 2683
rect -46 2611 -30 2645
rect 4 2611 20 2645
rect 646 2611 662 2645
rect 696 2611 712 2645
rect -30 2564 4 2611
rect 662 2566 696 2611
rect -46 1917 -30 1951
rect 4 1917 20 1951
rect 646 1917 662 1951
rect 696 1917 712 1951
rect -30 1870 4 1917
rect 662 1870 696 1917
rect -30 729 4 776
rect 662 729 696 776
rect -46 695 -30 729
rect 4 695 20 729
rect 646 695 662 729
rect 696 695 712 729
rect -30 35 4 82
rect 662 35 696 82
rect -46 1 -30 35
rect 4 1 20 35
rect 646 1 662 35
rect 696 1 712 35
rect -130 -37 -96 -11
rect 762 -37 796 -11
rect -130 -71 -70 -37
rect 736 -71 796 -37
<< viali >>
rect 662 2683 696 2717
rect -30 2611 4 2645
rect 662 2611 696 2645
rect -30 1917 4 1951
rect 662 1917 696 1951
rect -30 695 4 729
rect 662 695 696 729
rect -30 1 4 35
rect 662 1 696 35
rect -30 -71 4 -37
<< metal1 >>
rect 650 2717 708 2723
rect 650 2683 662 2717
rect 696 2683 708 2717
rect -42 2645 16 2651
rect -42 2611 -30 2645
rect 4 2611 16 2645
rect -42 2605 16 2611
rect 650 2645 708 2683
rect 650 2611 662 2645
rect 696 2611 708 2645
rect 650 2605 708 2611
rect -36 2564 10 2605
rect 656 2564 702 2605
rect -36 2552 97 2564
rect -49 2176 -39 2552
rect 13 2176 97 2552
rect -36 2164 97 2176
rect 310 2123 356 2564
rect 560 2557 702 2564
rect 560 2164 693 2557
rect 568 2123 614 2164
rect 310 2077 411 2123
rect 522 2077 614 2123
rect -42 1951 16 1957
rect -42 1917 -30 1951
rect 4 1917 16 1951
rect -42 1911 16 1917
rect -36 1870 10 1911
rect -36 1858 97 1870
rect -36 1482 49 1858
rect 101 1482 111 1858
rect -36 1470 97 1482
rect 52 1217 145 1263
rect 52 1176 97 1217
rect -36 776 97 1176
rect -36 735 10 776
rect -42 729 16 735
rect -42 695 -30 729
rect 4 695 16 729
rect -42 689 16 695
rect 310 569 356 2077
rect 650 1951 708 1957
rect 650 1917 662 1951
rect 696 1917 708 1951
rect 650 1911 708 1917
rect 656 1870 702 1911
rect 568 1470 701 1870
rect 568 1429 614 1470
rect 526 1383 614 1429
rect 568 1164 701 1176
rect 555 788 565 1164
rect 617 788 701 1164
rect 568 776 701 788
rect 656 735 702 776
rect 650 729 708 735
rect 650 695 662 729
rect 696 695 708 729
rect 650 689 708 695
rect 52 523 147 569
rect 264 523 356 569
rect 52 482 97 523
rect -36 82 97 482
rect 310 82 356 523
rect 568 470 701 482
rect 568 94 653 470
rect 705 94 715 470
rect 568 82 701 94
rect -36 41 10 82
rect 656 41 702 82
rect -42 35 16 41
rect -42 1 -30 35
rect 4 1 16 35
rect -42 -37 16 1
rect 650 35 708 41
rect 650 1 662 35
rect 696 1 708 35
rect 650 -5 708 1
rect -42 -71 -30 -37
rect 4 -71 16 -37
rect -42 -77 16 -71
<< via1 >>
rect -39 2176 13 2552
rect 49 1482 101 1858
rect 565 788 617 1164
rect 653 94 705 470
<< metal2 >>
rect -39 2552 13 2562
rect -39 2055 13 2176
rect -42 2046 14 2055
rect -42 1981 14 1990
rect 649 2048 709 2057
rect -39 658 13 1981
rect 649 1979 709 1988
rect 49 1858 101 1868
rect 49 1350 101 1482
rect 49 1298 617 1350
rect 565 1164 617 1298
rect 565 778 617 788
rect 653 665 705 1979
rect -52 598 -43 658
rect 17 598 26 658
rect 652 656 708 665
rect 652 591 708 600
rect 653 470 705 591
rect 653 84 705 94
<< via2 >>
rect -42 1990 14 2046
rect 649 1988 709 2048
rect -43 598 17 658
rect 652 600 708 656
<< metal3 >>
rect -47 2048 19 2051
rect 644 2048 714 2053
rect -47 2046 649 2048
rect -47 1990 -42 2046
rect 14 1990 649 2046
rect -47 1988 649 1990
rect 709 1988 714 2048
rect -47 1985 19 1988
rect 644 1983 714 1988
rect -48 658 22 663
rect 647 658 713 661
rect -48 598 -43 658
rect 17 656 713 658
rect 17 600 652 656
rect 708 600 713 656
rect 17 598 713 600
rect -48 593 22 598
rect 647 595 713 598
use sky130_fd_pr__pfet_01v8_2ZH9AN  sky130_fd_pr__pfet_01v8_2ZH9AN_0
timestamp 1729216653
transform 1 0 31 0 1 1670
box -109 -262 109 262
use sky130_fd_pr__pfet_01v8_2ZH9AN  sky130_fd_pr__pfet_01v8_2ZH9AN_1
timestamp 1729216653
transform 1 0 31 0 1 282
box -109 -262 109 262
use sky130_fd_pr__pfet_01v8_2ZH9AN  sky130_fd_pr__pfet_01v8_2ZH9AN_2
timestamp 1729216653
transform 1 0 635 0 1 282
box -109 -262 109 262
use sky130_fd_pr__pfet_01v8_2ZH9AN  sky130_fd_pr__pfet_01v8_2ZH9AN_3
timestamp 1729216653
transform 1 0 635 0 1 976
box -109 -262 109 262
use sky130_fd_pr__pfet_01v8_2ZH9AN  sky130_fd_pr__pfet_01v8_2ZH9AN_4
timestamp 1729216653
transform 1 0 31 0 1 976
box -109 -262 109 262
use sky130_fd_pr__pfet_01v8_2ZH9AN  sky130_fd_pr__pfet_01v8_2ZH9AN_5
timestamp 1729216653
transform 1 0 635 0 1 1670
box -109 -262 109 262
use sky130_fd_pr__pfet_01v8_2ZH9AN  sky130_fd_pr__pfet_01v8_2ZH9AN_6
timestamp 1729216653
transform 1 0 635 0 1 2364
box -109 -262 109 262
use sky130_fd_pr__pfet_01v8_2ZH9AN  sky130_fd_pr__pfet_01v8_2ZH9AN_7
timestamp 1729216653
transform 1 0 31 0 1 2364
box -109 -262 109 262
use sky130_fd_pr__pfet_01v8_SDE6B7  sky130_fd_pr__pfet_01v8_SDE6B7_0
timestamp 1729220975
transform 1 0 333 0 1 2364
box -323 -300 323 300
use sky130_fd_pr__pfet_01v8_SDE6B7  sky130_fd_pr__pfet_01v8_SDE6B7_1
timestamp 1729220975
transform 1 0 333 0 1 1670
box -323 -300 323 300
use sky130_fd_pr__pfet_01v8_SDE6B7  sky130_fd_pr__pfet_01v8_SDE6B7_2
timestamp 1729220975
transform 1 0 333 0 1 976
box -323 -300 323 300
use sky130_fd_pr__pfet_01v8_SDE6B7  sky130_fd_pr__pfet_01v8_SDE6B7_3
timestamp 1729220975
transform 1 0 333 0 1 282
box -323 -300 323 300
<< labels >>
flabel metal2 76 1394 76 1394 0 FreeSans 320 0 0 0 D1
port 0 nsew
flabel metal1 590 1416 590 1416 0 FreeSans 320 0 0 0 D2
port 1 nsew
flabel metal2 676 1364 676 1364 0 FreeSans 320 0 0 0 D5
port 2 nsew
flabel metal1 678 2670 678 2670 0 FreeSans 320 0 0 0 VDD
port 3 nsew
<< end >>
